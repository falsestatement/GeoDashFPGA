//-------------------------------------------------------------------------
//                                                                       --
//                                                                       --
//      For use with ECE 385 Lab 62                                       --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------


module lab62 (

      ///////// Clocks /////////
      input     MAX10_CLK1_50, 

      ///////// KEY /////////
      input    [ 1: 0]   KEY,

      ///////// SW /////////
      input    [ 9: 0]   SW,

      ///////// LEDR /////////
      output   [ 9: 0]   LEDR,

      ///////// HEX /////////
      output   [ 7: 0]   HEX0,
      output   [ 7: 0]   HEX1,
      output   [ 7: 0]   HEX2,
      output   [ 7: 0]   HEX3,
      output   [ 7: 0]   HEX4,
      output   [ 7: 0]   HEX5,

      ///////// SDRAM /////////
      output             DRAM_CLK,
      output             DRAM_CKE,
      output   [12: 0]   DRAM_ADDR,
      output   [ 1: 0]   DRAM_BA,
      inout    [15: 0]   DRAM_DQ,
      output             DRAM_LDQM,
      output             DRAM_UDQM,
      output             DRAM_CS_N,
      output             DRAM_WE_N,
      output             DRAM_CAS_N,
      output             DRAM_RAS_N,

      ///////// VGA /////////
      output             VGA_HS,
      output             VGA_VS,
      output   [ 3: 0]   VGA_R,
      output   [ 3: 0]   VGA_G,
      output   [ 3: 0]   VGA_B,


      ///////// ARDUINO /////////
      inout    [15: 0]   ARDUINO_IO,
      inout              ARDUINO_RESET_N 

);




logic Reset_h, vssig, blank, sync, VGA_Clk;


//=======================================================
//  REG/WIRE declarations
//=======================================================
	logic SPI0_CS_N, SPI0_SCLK, SPI0_MISO, SPI0_MOSI, USB_GPX, USB_IRQ, USB_RST, I2C_SDA_IN, I2C_SCL_IN, I2C_SDA_OE, I2C_SCL_OE;
	logic [3:0] hex_num_4, hex_num_3, hex_num_1, hex_num_0; //4 bit input hex digits
	logic [1:0] signs;
	logic [1:0] hundreds;
	logic [9:0] drawxsig, drawysig, ballxsig, ballysig, ballsizesig;
	logic [7:0] Red, Blue, Green;
	logic [7:0] keycode;
	logic [1:0] aud_mclk_ctr;

//=======================================================
//  Structural coding
//=======================================================
	assign ARDUINO_IO[10] = SPI0_CS_N;
	assign ARDUINO_IO[13] = SPI0_SCLK;
	assign ARDUINO_IO[11] = SPI0_MOSI;
	assign ARDUINO_IO[12] = 1'bZ;
	assign SPI0_MISO = ARDUINO_IO[12];
	
	assign ARDUINO_IO[9] = 1'bZ; 
	assign USB_IRQ = ARDUINO_IO[9];
		
	//Assignments specific to Circuits At Home UHS_20
	assign ARDUINO_RESET_N = USB_RST;
	assign ARDUINO_IO[7] = USB_RST;//USB reset 
	assign ARDUINO_IO[8] = 1'bZ; //this is GPX (set to input)
	assign USB_GPX = 1'b0;//GPX is not needed for standard USB host - set to 0 to prevent interrupt
	
	//Assign uSD CS to '1' to prevent uSD card from interfering with USB Host (if uSD card is plugged in)
	assign ARDUINO_IO[6] = 1'b1;
	
	//HEX drivers to convert numbers to HEX output
	HexDriver hex_driver4 (hex_num_4, HEX4[6:0]);
	assign HEX4[7] = 1'b1;
	
	HexDriver hex_driver3 (hex_num_3, HEX3[6:0]);
	assign HEX3[7] = 1'b1;
	
	HexDriver hex_driver1 (hex_num_1, HEX1[6:0]);
	assign HEX1[7] = 1'b1;
	
	HexDriver hex_driver0 (hex_num_0, HEX0[6:0]);
	assign HEX0[7] = 1'b1;
	
	//fill in the hundreds digit as well as the negative sign
	assign HEX5 = {1'b1, ~signs[1], 3'b111, ~hundreds[1], ~hundreds[1], 1'b1};
	assign HEX2 = {1'b1, ~signs[0], 3'b111, ~hundreds[0], ~hundreds[0], 1'b1};
	
	
	//Assign one button to reset
	assign {Reset_h}=~ (KEY[0]);

	//Our A/D converter is only 12 bit
	assign VGA_R = Red[7:4];
	assign VGA_B = Blue[7:4];
	assign VGA_G = Green[7:4];
	
	//I2C assignment stuff
	assign I2C_SDA_IN = ARDUINO_IO[14];
	assign I2C_SCL_IN = ARDUINO_IO[15];
	assign ARDUINO_IO[14] = I2C_SDA_OE ? 1'b0 : 1'bz;
	assign ARDUINO_IO[15] = I2C_SCL_OE ? 1'b0 : 1'bz;
	assign ARDUINO_IO[1] = 1'bz;
//	assign ARDUINO_IO[2] = ARDUINO_IO[1];
	
	//generate MCLK for SGTL5000
	assign ARDUINO_IO[3] = aud_mclk_ctr[1];
	always_ff @(posedge MAX10_CLK1_50) begin
		aud_mclk_ctr <= aud_mclk_ctr + 1;
	end
	
	logic[1:0] PLAYPLEASE;
	
	always_ff @ (posedge MAX10_CLK1_50)
	begin
		if(keycode == 8'h2c)
			PLAYPLEASE <= 2'b01;
		else 	if(collided)
			PLAYPLEASE <= 2'b10;
		else
			PLAYPLEASE <= 0;
	end

	
	
	lab62_soc u0 (
		.clk_clk                           (MAX10_CLK1_50),  //clk.clk
		.reset_reset_n                     (1'b1),           //reset.reset_n
		.altpll_0_locked_conduit_export    (),               //altpll_0_locked_conduit.export
		.altpll_0_phasedone_conduit_export (),               //altpll_0_phasedone_conduit.export
		.altpll_0_areset_conduit_export    (),               //altpll_0_areset_conduit.export
		.key_external_connection_export    (KEY),            //key_external_connection.export

		//SDRAM
		.sdram_clk_clk(DRAM_CLK),                            //clk_sdram.clk
		.sdram_wire_addr(DRAM_ADDR),                         //sdram_wire.addr
		.sdram_wire_ba(DRAM_BA),                             //.ba
		.sdram_wire_cas_n(DRAM_CAS_N),                       //.cas_n
		.sdram_wire_cke(DRAM_CKE),                           //.cke
		.sdram_wire_cs_n(DRAM_CS_N),                         //.cs_n
		.sdram_wire_dq(DRAM_DQ),                             //.dq
		.sdram_wire_dqm({DRAM_UDQM,DRAM_LDQM}),              //.dqm
		.sdram_wire_ras_n(DRAM_RAS_N),                       //.ras_n
		.sdram_wire_we_n(DRAM_WE_N),                         //.we_n

		//USB SPI	
		.spi0_SS_n(SPI0_CS_N),
		.spi0_MOSI(SPI0_MOSI),
		.spi0_MISO(SPI0_MISO),
		.spi0_SCLK(SPI0_SCLK),
		
		//USB GPIO
		.usb_rst_export(USB_RST),
		.usb_irq_export(USB_IRQ),
		.usb_gpx_export(USB_GPX),
		
		//LEDs and HEX
		.hex_digits_export({hex_num_4, hex_num_3, hex_num_1, hex_num_0}),
		.leds_export({hundreds, signs, LEDR}),
		.keycode_export(keycode),
		
		//i2c stuff
		.i2c_serial_out_sda_in(I2C_SDA_IN),          //          i2c_serial_out.sda_in
		.i2c_serial_out_scl_in(I2C_SCL_IN),          //                        .scl_in
		.i2c_serial_out_sda_oe(I2C_SDA_OE),          //                        .sda_oe
		.i2c_serial_out_scl_oe(I2C_SCL_OE)
	 );


I2S_Interface i2s(
	 .PLAYPLEASE(PLAYPLEASE),
    .LRCLK(ARDUINO_IO[4]), .SCLK(ARDUINO_IO[5]),
    .D_OUT(ARDUINO_IO[2])
	 );
	 
//instantiate a vga_controller, ball, and color_mapper here with the ports

vga_controller vga( .Clk(MAX10_CLK1_50),
										 .Reset(Reset_h),
										 //output logic
										 .hs(VGA_HS),
										 .vs(VGA_VS),
										 .pixel_clk(VGA_Clk),
										 .blank(blank),
										 .sync(sync),
										 //outputs
										 .DrawX(drawxsig),
										 .DrawY(drawysig)
										);

color_mapper cmap( 					.BallX(ballxsig),
									.BallY(ballysig),
									.Triangle_X(trianglexsig),
									.Triangle_Y(triangleysig),
									.Column_X(columnxsig),
									.DrawX(drawxsig),
									.DrawY(drawysig),
									.is_flipped(is_flipped),
									.will_collide(will_collide),
									.Ball_size(ballsizesig),
									//outputs
									.Red(Red),
									.Green(Green),
									.Blue(Blue)
								 );
								 
ball ball_obj( .Reset(Reset_h),
			   .frame_clk(VGA_VS),
				.keycode(keycode),
				.game(game_state),
				.collided(collided),
				.startRandom(startRandom),
				//outputs
				.BallX(ballxsig),
				.BallY(ballysig),
				.BallS(ballsizesig)
			 );


logic is_flipped, collided, colTri1, colColumn;
logic [1:0] game_state;
logic [10:0] trianglexsig, triangleysig, columnxsig;

assign collided = colTri1 || colColumn;
// assign columnxsig = 310;
// assign trianglexsig = 500;
// assign triangleysig = 317;

logic [26:0] random_clk_ctr;
//logic [4:0] random_number;

logic startRandom, spT1, spC;

// fibonacci_lfsr randGen (
//   .clk (MAX10_CLK1_50),
//   .rst_n (Reset_h),
//   .data (random_number)
// );
//
//initial begin
//	random_number = 23;
//end

always_ff @(posedge MAX10_CLK1_50) begin
		random_clk_ctr <= random_clk_ctr + 1;
//		random_number = next_item(random_number);
	end


logic [2:0] PathStep;
always_ff @ (posedge random_clk_ctr[24])
begin
	if(startRandom) begin
		unique case (PathStep)
			0:
			begin
				if(trianglexsig == 640 && columnxsig == 640 && !collided) begin
					spT1 <= 1;
					PathStep <= PathStep + 1;
				end
				else begin
					spT1 <= 0;
					spC <= 0;
				end
			end
			1:
			begin
				if(trianglexsig == 640 && columnxsig == 640 && !collided) begin
					spT1 <= 1;
					PathStep <= PathStep + 1;
				end
				else begin
					spT1 <= 0;
					spC <= 0;
				end
			end
			2:
			begin
				if(trianglexsig == 640 && columnxsig == 640 && !collided) begin
					spC <= 1;
					PathStep <= PathStep + 1;
				end
				else begin
					spT1 <= 0;
					spC <= 0;
				end
			end
			3:
			begin
				if(trianglexsig == 640 && columnxsig == 640 && !collided) begin
					spT1 <= 1;
					PathStep <= PathStep + 1;
				end
				else begin
					spT1 <= 0;
					spC <= 0;
				end
			end
			4:
			begin
				if(trianglexsig == 640 && columnxsig == 640 && !collided) begin
					spT1 <= 1;
					PathStep <= PathStep + 1;
				end
				else begin
					spT1 <= 0;
					spC <= 0;
				end
			end
			5:
			begin
				if(trianglexsig == 640 && columnxsig == 640 && !collided) begin
					spC <= 1;
					PathStep <= PathStep + 1;
				end
				else begin
					spT1 <= 0;
					spC <= 0;
				end
			end
			6:
			begin
				if(trianglexsig == 640 && columnxsig == 640 && !collided) begin
					spT1 <= 1;
					PathStep <= PathStep + 1;
				end
				else begin
					spT1 <= 0;
					spC <= 0;
				end
			end
			7:
			begin
				if(trianglexsig == 640 && columnxsig == 640 && !collided) begin
					spT1 <= 1;
					PathStep <= PathStep + 1;
				end
				else begin
					spT1 <= 0;
					spC <= 0;
				end
			end
		endcase
	end
end

assign is_flipped = game_state[0];

obstacle_triangle triangle1(
    .is_flipped(is_flipped), 
	.start_moving(spT1),
    .Player_Y(ballysig), 
	.Player_size(ballsizesig),
    .Reset(Reset_h), 
	.frame_clk(VGA_VS),
	.Triangle_X(trianglexsig), 
	.Triangle_Y(triangleysig),
	.will_collide(colTri1)
);

obstacle_column flip_column
(
    .start_moving(spC),
    .game_state(game_state),
    .Player_Y(ballysig), 
	.Player_size(ballsizesig),
    .Reset(Reset_h), 
	.frame_clk(VGA_VS),
	.Column_X(columnxsig),
	.will_collide(colColumn), 
	.passed_through()
);

endmodule


// credit to https://stackoverflow.com/questions/67361956/how-to-generate-a-synthesizable-pseudo-random-generator-from-1-to-52-system-veri
function [5:0] next_item(input logic [5:0] v);
  if(v < 26) begin
    next_item = (v << 1); // 2 * v % 53 = 2 * v
  end
  else if(v > 26) begin
    // (2 * v) % 53 = (2 * v - 52 - 1) % 53 = 2 * (v - 26) - 1
    next_item = (((v - 26) << 2) - 1);
  end
  else begin
    // v = 26, you want to exclude 2 * v % 53 = 52, so we skip it
    // by applying the next item again, and it will be 
    next_item = 51;
  end
endfunction